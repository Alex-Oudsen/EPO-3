library IEEE;
use IEEE.std_logic_1164.ALL;

entity tb_compare is
end tb_compare;


