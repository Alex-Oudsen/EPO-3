library IEEE;
use IEEE.std_logic_1164.ALL;

entity ram_tb is
end ram_tb;


