library IEEE;
use IEEE.std_logic_1164.ALL;

entity controller_tb is
end controller_tb;
