-- Alex Oudsen, 4325494

library ieee;
use ieee.std_logic_1164.all;

entity mod24_tel_tb is
end mod24_tel_tb;
