library IEEE;
use IEEE.std_logic_1164.ALL;

entity top_top_tb is
end top_top_tb;
