configuration fifo_behaviour_cfg of fifo is
   for behaviour
   end for;
end fifo_behaviour_cfg;


