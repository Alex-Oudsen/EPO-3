library IEEE;
use IEEE.std_logic_1164.ALL;

entity dcf_lcd_tb is
end dcf_lcd_tb;


