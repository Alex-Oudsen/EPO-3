-- Alex Oudsen, 4325494

library ieee;
use ieee.std_logic_1164.all;

entity autosyncklok_tb is
end entity autosyncklok_tb;