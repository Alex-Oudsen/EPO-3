library IEEE;
use IEEE.std_logic_1164.ALL;

entity licht_tb is
end licht_tb;


