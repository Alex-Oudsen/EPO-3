configuration ram_behaviour_cfg of ram is
   for behaviour
   end for;
end ram_behaviour_cfg;


