library IEEE;
use IEEE.std_logic_1164.ALL;

entity wektijd_tb is
end wektijd_tb;


