library IEEE;
use IEEE.std_logic_1164.ALL;

entity tijd_tb is
end tijd_tb;


