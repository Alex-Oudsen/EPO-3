-- Alex Oudsen, 4325494

library ieee;
use ieee.std_logic_1164.all;

entity parity_tb is
end parity_tb;