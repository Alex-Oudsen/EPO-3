library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of datum_tb is
begin
end behaviour;


