configuration send_cntrl_tb_behaviour_cfg of send_cntrl_tb is
   for behaviour
   end for;
end send_cntrl_tb_behaviour_cfg;


