library IEEE;
use IEEE.std_logic_1164.ALL;

entity counter_tb is
end counter_tb;


