configuration send_bus_behaviour_cfg of send_bus is
   for behaviour
   end for;
end send_bus_behaviour_cfg;


