-- Alex Oudsen, 4325494

library ieee;
use ieee.std_logic_1164.all;

entity parity_check_tb is
end parity_check_tb;