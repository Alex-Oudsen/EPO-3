configuration send_control_behaviour_cfg of send_control is
   for behaviour
   end for;
end send_control_behaviour_cfg;


