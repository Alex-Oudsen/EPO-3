configuration send_bus_tb_behaviour_cfg of send_bus_tb is
   for behaviour
   end for;
end send_bus_tb_behaviour_cfg;


