library IEEE;
use IEEE.std_logic_1164.ALL;

entity tb_fifo_ctr is
end tb_fifo_ctr;


