-- Alex Oudsen, 4325494

library ieee;
use ieee.std_logic_1164.all;

entity bcd2bin_tb is
end bcd2bin_tb;