library IEEE;
use IEEE.std_logic_1164.ALL;

entity menu_scherm_tb is
end menu_scherm_tb;


