library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of controller is
signal wekdata_in, wekdata_out : std_logic_vector(13 downto 0);
begin
end behaviour;


