-- Alex Oudsen, 4325494

library ieee;
use ieee.std_logic_1164.all;

entity dcf77_tb is
end dcf77_tb;