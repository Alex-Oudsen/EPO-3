library IEEE;
use IEEE.std_logic_1164.ALL;

entity lcd_top_tb is
end lcd_top_tb;
