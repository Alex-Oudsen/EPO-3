-- Alex Oudsen, 4325494

library ieee;
use ieee.std_logic_1164.all;

entity klokdeler_tb is
end entity klokdeler_tb;