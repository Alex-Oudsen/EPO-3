library ieee;

entity alu_tb is
end entity alu_tb;
