configuration tijd_behaviour_cfg of tijd is
   for behaviour
   end for;
end tijd_behaviour_cfg;


