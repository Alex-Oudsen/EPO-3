-- Alex Oudsen, 4325494

library ieee;
use ieee.std_logic_1164.all;

entity dcf_counter_tb is
end dcf_counter_tb;
