-- Alex Oudsen, 4325494

library ieee;
use ieee.std_logic_1164.all;

entity edge_detect_tb is
end entity edge_detect_tb;