library ieee;
use ieee.std_logic_1164.all;

entity alu_tb is
end entity alu_tb;

