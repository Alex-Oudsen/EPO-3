library IEEE;
use IEEE.std_logic_1164.ALL;

entity send_cntrl_tb is
end send_cntrl_tb;


