configuration fifo_synthesised_cfg of fifo is
   for synthesised
   end for;
end fifo_synthesised_cfg;


