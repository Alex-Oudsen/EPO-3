library IEEE;
use IEEE.std_logic_1164.ALL;

entity datum_tb is
end datum_tb;


