configuration fifo_totaal_extracted_cfg of fifo_totaal is
   for extracted
   end for;
end fifo_totaal_extracted_cfg;


