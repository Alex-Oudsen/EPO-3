-- Alex Oudsen, 4325494

library ieee;
use ieee.std_logic_1164.all;

entity synctime_tb is
end synctime_tb;
