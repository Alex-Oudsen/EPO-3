library IEEE;
use IEEE.std_logic_1164.ALL;

entity send_bus_tb is
end send_bus_tb;


