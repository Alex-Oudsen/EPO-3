library ieee;
use ieee.std_logic_1164.all;

entity wake_up_tb is
end wake_up_tb;


