library IEEE;
use IEEE.std_logic_1164.ALL;

entity alarm is
   port(clk       :in    std_logic;
        reset     :in    std_logic;
        sec       :in    std_logic;
        licht     :in    std_logic;
        pwm_signal:out   std_logic);
end alarm;


