configuration send_bus_synthesised_cfg of send_bus is
   for synthesised
   end for;
end send_bus_synthesised_cfg;


