library IEEE;
use IEEE.std_logic_1164.ALL;

entity tb_alarm is
end tb_alarm;


