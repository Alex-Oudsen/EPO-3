library IEEE;
use IEEE.std_logic_1164.ALL;

entity pwm_tb is
end pwm_tb;


