library IEEE;
use IEEE.std_logic_1164.ALL;

entity geluid_tb is
end geluid_tb;


