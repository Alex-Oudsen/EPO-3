library IEEE;
use IEEE.std_logic_1164.ALL;

entity totaal_tb is
end totaal_tb;


